module top(
    input i_clk,
    input i_clk_1Hz,
    output [6:0] o_hex,
);



7_segment_display 7_segment_display_Inst
(.i_3bit_bin_num(r_num),


)
